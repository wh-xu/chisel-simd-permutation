../generated/simd_permutation_network.sv