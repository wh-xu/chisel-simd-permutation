../generated/SimdPermutation.sv